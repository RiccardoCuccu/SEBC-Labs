library ieee ;
  use ieee.std_logic_1164.all ;
  use ieee.numeric_std.all ;

package constants is
   constant N_BIT : integer := 32;
end constants;
